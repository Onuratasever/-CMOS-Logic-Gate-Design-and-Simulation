magic
tech scmos
timestamp 1730402689
<< nwell >>
rect -15 -7 17 18
<< ntransistor >>
rect -4 -77 -2 -73
rect 2 -77 4 -73
<< ptransistor >>
rect -4 -1 -2 7
rect 4 -1 6 7
<< ndiffusion >>
rect -5 -77 -4 -73
rect -2 -77 2 -73
rect 4 -77 5 -73
<< pdiffusion >>
rect -5 -1 -4 7
rect -2 -1 -1 7
rect 3 -1 4 7
rect 6 -1 7 7
<< ndcontact >>
rect -9 -77 -5 -73
rect 5 -77 9 -73
<< pdcontact >>
rect -9 -1 -5 7
rect -1 -1 3 7
rect 7 -1 11 7
<< psubstratepcontact >>
rect -9 -85 -5 -81
rect 5 -85 9 -81
<< nsubstratencontact >>
rect -9 11 -5 15
rect 7 11 11 15
<< polysilicon >>
rect -4 7 -2 10
rect 4 7 6 10
rect -4 -73 -2 -1
rect 4 -70 6 -1
rect 2 -72 6 -70
rect 2 -73 4 -72
rect -4 -80 -2 -77
rect 2 -80 4 -77
<< polycontact >>
rect -8 -18 -4 -14
rect 6 -12 10 -8
<< metal1 >>
rect -5 11 7 15
rect -9 7 -5 11
rect 7 7 11 11
rect -1 -16 3 -1
rect -1 -20 9 -16
rect 5 -57 9 -20
rect 5 -61 11 -57
rect 5 -73 9 -61
rect -9 -81 -5 -77
rect -5 -85 5 -81
<< labels >>
rlabel metal1 0 -83 0 -83 1 gnd
rlabel polycontact -6 -16 -6 -16 1 input1
rlabel polycontact 8 -10 8 -10 1 input2
rlabel metal1 1 13 1 13 5 vddd
rlabel metal1 9 -59 9 -59 1 output
<< end >>
