magic
tech scmos
timestamp 1730406563
<< nwell >>
rect -7 -11 17 14
<< ntransistor >>
rect 4 -81 6 -77
<< ptransistor >>
rect 4 -5 6 3
<< ndiffusion >>
rect 3 -81 4 -77
rect 6 -81 7 -77
<< pdiffusion >>
rect 3 -5 4 3
rect 6 -5 7 3
<< ndcontact >>
rect -1 -81 3 -77
rect 7 -81 11 -77
<< pdcontact >>
rect -1 -5 3 3
rect 7 -5 11 3
<< psubstratepcontact >>
rect -1 -89 3 -85
rect 7 -89 11 -85
<< nsubstratencontact >>
rect -1 7 3 11
rect 7 7 11 11
<< polysilicon >>
rect 4 3 6 6
rect 4 -77 6 -5
rect 4 -84 6 -81
<< polycontact >>
rect 0 -17 4 -13
<< metal1 >>
rect 3 7 7 11
rect -1 3 3 7
rect 7 -14 11 -5
rect 7 -18 13 -14
rect 7 -77 11 -18
rect -1 -85 3 -81
rect 3 -89 7 -85
<< labels >>
rlabel polycontact 2 -15 2 -15 1 input
rlabel metal1 10 -16 10 -16 1 output
rlabel metal1 5 9 5 9 5 vddd
rlabel metal1 5 -87 5 -87 1 gnd
<< end >>
